module datapath ()

endmodule