module PS2_Decoder ()

    


endmodule 

