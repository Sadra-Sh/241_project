module control ()

endmodule

module datapath ()

endmodule