module datapath(
    input clk,
    input Reset,
    input [7:0] data_in,
    input ld_alu_out,
    input ld_x, ld_a, ld_b, ld_c,
    input ld_r,
    input alu_op,
    input [1:0] alu_select_a, alu_select_b,
    output reg [7:0] data_result
    );
    // input registers
    reg [7:0] a, b, c, x;
    // output of the alu
    reg [7:0] alu_out;
    // alu input muxes
    reg [7:0] alu_a, alu_b;
    // Registers a, b, c, x with respective input logic
    always@(posedge clk) begin
    if(Reset) begin
    a <= 8'b0;
    b <= 8'b0;
    c <= 8'b0;
    x <= 8'b0;
    end
    else begin
    if(ld_a)
    a <= ld_alu_out ? alu_out : data_in; // load alu_out if
    load_alu_out signal is high, otherwise load from data_in
    if(ld_b)
    b <= ld_alu_out ? alu_out : data_in; // load alu_out if
    load_alu_out signal is high, otherwise load from data_in
    if(ld_x)
    x <= data_in;
    if(ld_c)
    c <= data_in;
    end
    end
    // Output result register
    always@(posedge clk) begin
    if(Reset) begin
    data_result <= 8'b0;
    end
    else
    if(ld_r)
    data_result <= alu_out;
    end
    // The ALU input multiplexers
    always @(*)
    begin
    case (alu_select_a)
    2'd0:
    alu_a = a;
    2'd1:
    alu_a = b;
    2'd2:
    alu_a = c;
    2'd3:
    alu_a = x;
    default: alu_a = 8'b0;
    endcase
    case (alu_select_b)
    2'd0:
    alu_b = a;
    2'd1:
    alu_b = b;
    2'd2:
    alu_b = c;
    2'd3:
    alu_b = x;
    default: alu_b = 8'b0;
    endcase
    end
    // The ALU
    always @(*)
    begin : ALU
    // alu
    case (alu_op)
    0: begin
    alu_out = alu_a + alu_b; //performs addition
    end
    1: begin
    alu_out = alu_a * alu_b; //performs multiplication
    end
    default: alu_out = 8'b0;
    endcase
    end
endmodule
